module gi

#flag `pkg-config --cflags gobject-introspection-1.0` `pkg-config --libs gobject-introspection-1.0`

#include <girepository.h>
