module gi
