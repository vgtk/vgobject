module gi

pub struct CallbackInfo {
	c &GICallbackInfo
}
