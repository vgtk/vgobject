module gi

type gi__ConstantInfo BaseInfo

// TODO
